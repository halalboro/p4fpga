`timescale 1ns / 1ps

// =============================================================================
// QoS (Quality of Service) Testbench
//
// Tests DSCP marking based on IP protocol (qos.p4):
// - LPM match on IPv4 destination address
// - Conditional QoS marking:
//   - UDP (protocol=17) -> Expedited Forwarding (diffserv=46)
//   - TCP (protocol=6)  -> Voice Admit (diffserv=44)
// - Actions: ipv4_forward, drop, NoAction
// =============================================================================

module tb_user;
    // ==========================================
    // Clock and Reset
    // ==========================================
    logic aclk = 1'b1;
    logic aresetn = 1'b0;

    localparam CLK_PERIOD = 4ns;  // 250 MHz
    always #(CLK_PERIOD/2) aclk = ~aclk;

    initial begin
        aresetn = 1'b0;
        #100ns aresetn = 1'b1;
    end

    // ==========================================
    // Parameters
    // ==========================================
    localparam DATA_WIDTH = 512;
    localparam KEEP_WIDTH = DATA_WIDTH/8;
    localparam ACTION_DATA_WIDTH = 128;

    // Protocol constants
    localparam [7:0] PROTO_ICMP = 8'd1;
    localparam [7:0] PROTO_TCP  = 8'd6;
    localparam [7:0] PROTO_UDP  = 8'd17;

    // Expected DSCP values
    localparam [5:0] DSCP_DEFAULT = 6'd0;
    localparam [5:0] DSCP_EF      = 6'd46;  // Expedited Forwarding (UDP)
    localparam [5:0] DSCP_VA      = 6'd44;  // Voice Admit (TCP)

    // ==========================================
    // AXI-Stream interfaces
    // ==========================================
    logic [DATA_WIDTH-1:0]   s_axis_tdata;
    logic [KEEP_WIDTH-1:0]   s_axis_tkeep;
    logic                    s_axis_tvalid;
    logic                    s_axis_tlast;
    logic                    s_axis_tready;

    logic [DATA_WIDTH-1:0]   m_axis_tdata;
    logic [KEEP_WIDTH-1:0]   m_axis_tkeep;
    logic                    m_axis_tvalid;
    logic                    m_axis_tlast;
    logic                    m_axis_tready;

    // ==========================================
    // Table programming signals
    // ==========================================
    logic        table_wr_en;
    logic [9:0]  table_wr_addr;
    logic        table_entry_valid;
    logic [31:0] table_entry_prefix;
    logic [5:0]  table_entry_prefix_len;
    logic [2:0]  table_entry_action;
    logic [ACTION_DATA_WIDTH-1:0] table_entry_action_data;

    // Ingress port
    logic [8:0]  ingress_port;

    // ==========================================
    // Statistics
    // ==========================================
    logic [31:0] packet_count, dropped_count, forwarded_count;
    logic        pipeline_drop;

    int packets_sent = 0;
    int packets_received = 0;

    // ==========================================
    // Parser output signals
    // ==========================================
    logic        ethernet_valid;
    logic [47:0] eth_dst_addr, eth_src_addr;
    logic [15:0] eth_type;
    logic        ipv4_valid, tcp_valid, udp_valid;
    logic [3:0]  ipv4_version, ipv4_ihl;
    logic [5:0]  ipv4_diffserv;
    logic [1:0]  ipv4_ecn;
    logic [15:0] ipv4_totalLen, ipv4_identification;
    logic [2:0]  ipv4_flags;
    logic [12:0] ipv4_fragOffset;
    logic [7:0]  ipv4_ttl, ipv4_protocol;
    logic [15:0] ipv4_hdrChecksum;
    logic [31:0] ipv4_src_addr, ipv4_dst_addr;
    logic [15:0] tcp_src_port, tcp_dst_port;
    logic [15:0] udp_src_port, udp_dst_port;

    logic [DATA_WIDTH-1:0]  parser_payload_data;
    logic [KEEP_WIDTH-1:0]  parser_payload_keep;
    logic                   parser_payload_valid, parser_payload_last, parser_payload_ready;
    logic [15:0]            parser_packet_length;
    logic [8:0]             parser_ingress_port;

    // ==========================================
    // Pipeline signals
    // ==========================================
    logic [DATA_WIDTH-1:0]  pipeline_data;
    logic [KEEP_WIDTH-1:0]  pipeline_keep;
    logic                   pipeline_last, pipeline_valid, pipeline_ready;
    logic [8:0]             pipeline_egress_port, pipeline_egress_port_d;
    logic                   pipeline_header_modified;
    logic [5:0]             pipeline_ipv4_diffserv;
    logic [1:0]             pipeline_ipv4_ecn;
    logic [7:0]             pipeline_ipv4_ttl;
    logic [47:0]            pipeline_eth_dst, pipeline_eth_src;

    // ==========================================
    // Action IDs (from P4 program)
    // ==========================================
    localparam ACTION_FORWARD  = 3'd0;   // ipv4_forward
    localparam ACTION_DROP     = 3'd1;   // drop
    localparam ACTION_NOACTION = 3'd2;   // NoAction
    // Conditional actions generated by compiler
    localparam ACTION_EF       = 3'd14;  // expedited_forwarding (UDP)
    localparam ACTION_VA       = 3'd16;  // voice_admit (TCP) - Note: truncated to 3 bits

    // ==========================================
    // Parser Instance
    // ==========================================
    parser #(
        .DATA_WIDTH(DATA_WIDTH),
        .PARSER_CONFIG(8'b00100101)  // Ethernet + IPv4 + UDP
    ) parser_inst (
        .aclk(aclk),
        .aresetn(aresetn),
        .s_axis_tdata(s_axis_tdata),
        .s_axis_tkeep(s_axis_tkeep),
        .s_axis_tvalid(s_axis_tvalid),
        .s_axis_tlast(s_axis_tlast),
        .s_axis_tready(s_axis_tready),
        .eth_dst_addr(eth_dst_addr),
        .eth_src_addr(eth_src_addr),
        .eth_ether_type(eth_type),
        .eth_valid(ethernet_valid),
        .vlan_pcp(),
        .vlan_dei(),
        .vlan_vid(),
        .vlan_ether_type(),
        .vlan_valid(),
        .ipv4_version(ipv4_version),
        .ipv4_ihl(ipv4_ihl),
        .ipv4_diffserv(ipv4_diffserv),
        .ipv4_ecn(ipv4_ecn),
        .ipv4_total_len(ipv4_totalLen),
        .ipv4_identification(ipv4_identification),
        .ipv4_flags(ipv4_flags),
        .ipv4_frag_offset(ipv4_fragOffset),
        .ipv4_ttl(ipv4_ttl),
        .ipv4_protocol(ipv4_protocol),
        .ipv4_hdr_checksum(ipv4_hdrChecksum),
        .ipv4_src_addr(ipv4_src_addr),
        .ipv4_dst_addr(ipv4_dst_addr),
        .ipv4_valid(ipv4_valid),
        .ipv6_version(),
        .ipv6_traffic_class(),
        .ipv6_flow_label(),
        .ipv6_payload_len(),
        .ipv6_next_hdr(),
        .ipv6_hop_limit(),
        .ipv6_src_addr(),
        .ipv6_dst_addr(),
        .ipv6_valid(),
        .tcp_src_port(tcp_src_port),
        .tcp_dst_port(tcp_dst_port),
        .tcp_seq_no(),
        .tcp_ack_no(),
        .tcp_data_offset(),
        .tcp_reserved(),
        .tcp_flags(),
        .tcp_window(),
        .tcp_checksum(),
        .tcp_urgent_ptr(),
        .tcp_valid(tcp_valid),
        .udp_src_port(udp_src_port),
        .udp_dst_port(udp_dst_port),
        .udp_length(),
        .udp_checksum(),
        .udp_valid(udp_valid),
        .vxlan_flags(),
        .vxlan_reserved(),
        .vxlan_vni(),
        .vxlan_reserved2(),
        .vxlan_valid(),
        .payload_data(parser_payload_data),
        .payload_keep(parser_payload_keep),
        .payload_valid(parser_payload_valid),
        .payload_last(parser_payload_last),
        .packet_length(parser_packet_length),
        .ingress_port(parser_ingress_port)
    );

    // Egress port delay for feedback
    always_ff @(posedge aclk) pipeline_egress_port_d <= pipeline_egress_port;

    // ==========================================
    // Match-Action Pipeline Instance
    // ==========================================
    match_action #(
        .DATA_WIDTH(DATA_WIDTH),
        .TABLE_SIZE(1024),
        .KEY_WIDTH(32),                // 32-bit IPv4 address for LPM
        .ACTION_DATA_WIDTH(ACTION_DATA_WIDTH),
        .ACTION_CONFIG(8'b01000111),   // Forward, Drop, Modify, SET_FIELD
        .EGRESS_CONFIG(8'b00000000),   // No special egress features
        .NUM_REGISTERS(1024)
    ) match_action_inst (
        .aclk(aclk),
        .aresetn(aresetn),
        .metadata_in(64'd0),
        .metadata_out(),
        .packet_in(parser_payload_data),
        .packet_keep_in(parser_payload_keep),
        .packet_last_in(parser_payload_last),
        .packet_valid_in(parser_payload_valid),
        .packet_ready_out(parser_payload_ready),
        .ingress_port_in(ingress_port),
        .ipv4_valid(ipv4_valid),
        .eth_dst_addr(eth_dst_addr),
        .eth_src_addr(eth_src_addr),
        .ipv4_ttl(ipv4_ttl),
        .ipv4_src_addr(ipv4_src_addr),
        .ipv4_dst_addr(ipv4_dst_addr),
        .ipv4_src_port(udp_src_port),
        .ipv4_dst_port(udp_dst_port),
        .ipv4_protocol(ipv4_protocol),
        .ipv4_diffserv(ipv4_diffserv),
        .ipv4_ecn(ipv4_ecn),
        .packet_length(parser_packet_length),
        .mcast_grp(),
        .enq_qdepth(19'd0),
        .egress_port_id(pipeline_egress_port_d),
        .packet_out(pipeline_data),
        .packet_keep_out(pipeline_keep),
        .packet_last_out(pipeline_last),
        .packet_valid_out(pipeline_valid),
        .packet_ready_in(pipeline_ready),
        .out_ipv4_diffserv(pipeline_ipv4_diffserv),
        .out_ipv4_ecn(pipeline_ipv4_ecn),
        .out_ipv4_ttl(pipeline_ipv4_ttl),
        .out_eth_dst_addr(pipeline_eth_dst),
        .out_eth_src_addr(pipeline_eth_src),
        .drop(pipeline_drop),
        .egress_port(pipeline_egress_port),
        .header_modified(pipeline_header_modified),
        .ecn_marked(),
        .table_write_enable(table_wr_en),
        .table_write_addr(table_wr_addr),
        .table_entry_valid(table_entry_valid),
        .table_entry_key(table_entry_prefix),
        .table_entry_prefix_len(table_entry_prefix_len),
        .table_entry_action(table_entry_action),
        .table_entry_action_data(table_entry_action_data),
        .packet_count(packet_count),
        .dropped_count(dropped_count),
        .forwarded_count(forwarded_count)
    );

    // ==========================================
    // Deparser Instance
    // ==========================================
    deparser #(
        .DATA_WIDTH(DATA_WIDTH),
        .DEPARSER_CONFIG(16'h0085)  // Ethernet + IPv4 + checksum update
    ) deparser_inst (
        .aclk(aclk),
        .aresetn(aresetn),
        .eth_dst_addr(pipeline_eth_dst),
        .eth_src_addr(pipeline_eth_src),
        .eth_ether_type(eth_type),
        .eth_valid(ethernet_valid),
        .vlan_pcp(3'b0),
        .vlan_dei(1'b0),
        .vlan_vid(12'b0),
        .vlan_ether_type(16'b0),
        .vlan_valid(1'b0),
        .ipv4_version(ipv4_version),
        .ipv4_ihl(ipv4_ihl),
        .ipv4_diffserv(pipeline_ipv4_diffserv),
        .ipv4_ecn(pipeline_ipv4_ecn),
        .ipv4_total_len(ipv4_totalLen),
        .ipv4_identification(ipv4_identification),
        .ipv4_flags(ipv4_flags),
        .ipv4_frag_offset(ipv4_fragOffset),
        .ipv4_ttl(pipeline_ipv4_ttl),
        .ipv4_protocol(ipv4_protocol),
        .ipv4_hdr_checksum(ipv4_hdrChecksum),
        .ipv4_src_addr(ipv4_src_addr),
        .ipv4_dst_addr(ipv4_dst_addr),
        .ipv4_valid(ipv4_valid),
        .ipv6_version(4'd0),
        .ipv6_traffic_class(8'd0),
        .ipv6_flow_label(20'd0),
        .ipv6_payload_len(16'd0),
        .ipv6_next_hdr(8'd0),
        .ipv6_hop_limit(8'd0),
        .ipv6_src_addr(128'd0),
        .ipv6_dst_addr(128'd0),
        .ipv6_valid(1'b0),
        .tcp_src_port(16'd0),
        .tcp_dst_port(16'd0),
        .tcp_seq_no(32'd0),
        .tcp_ack_no(32'd0),
        .tcp_data_offset(4'd5),
        .tcp_reserved(3'd0),
        .tcp_flags(9'd0),
        .tcp_window(16'd0),
        .tcp_checksum(16'd0),
        .tcp_urgent_ptr(16'd0),
        .tcp_valid(1'b0),
        .udp_src_port(16'd0),
        .udp_dst_port(16'd0),
        .udp_length(16'd0),
        .udp_checksum(16'd0),
        .udp_valid(1'b0),
        .vxlan_flags(8'd0),
        .vxlan_reserved(24'd0),
        .vxlan_vni(24'd0),
        .vxlan_reserved2(8'd0),
        .vxlan_valid(1'b0),
        .s_axis_tdata(pipeline_data),
        .s_axis_tkeep(pipeline_keep),
        .s_axis_tvalid(pipeline_valid),
        .s_axis_tlast(pipeline_last),
        .s_axis_tready(pipeline_ready),
        .drop_packet(pipeline_drop),
        .m_axis_tdata(m_axis_tdata),
        .m_axis_tkeep(m_axis_tkeep),
        .m_axis_tvalid(m_axis_tvalid),
        .m_axis_tlast(m_axis_tlast),
        .m_axis_tready(m_axis_tready)
    );

    // ==========================================
    // Byte swap functions
    // ==========================================
    function automatic [47:0] bswap48(input [47:0] val);
        bswap48 = {val[7:0], val[15:8], val[23:16], val[31:24], val[39:32], val[47:40]};
    endfunction

    function automatic [31:0] bswap32(input [31:0] val);
        bswap32 = {val[7:0], val[15:8], val[23:16], val[31:24]};
    endfunction

    function automatic [15:0] bswap16(input [15:0] val);
        bswap16 = {val[7:0], val[15:8]};
    endfunction

    // ==========================================
    // Task: Configure LPM route entry
    // ==========================================
    task configure_route(
        input [9:0]  addr,
        input [31:0] prefix,
        input [5:0]  prefix_len,
        input [2:0]  action_id,
        input [47:0] dst_mac,
        input [8:0]  egress_p
    );
        @(posedge aclk);
        table_wr_en            <= 1'b1;
        table_wr_addr          <= addr;
        table_entry_valid      <= 1'b1;
        table_entry_prefix     <= prefix;
        table_entry_prefix_len <= prefix_len;
        table_entry_action     <= action_id;
        // action_data format: [103:96]=egress_port, [47:0]=dst_mac
        table_entry_action_data <= {24'd0, egress_p[7:0], 48'd0, dst_mac};

        @(posedge aclk);
        table_wr_en <= 1'b0;
        @(posedge aclk);

        $display("[%0t] Route configured: addr=%0d prefix=%08h/%0d action=%0d port=%0d",
                 $time, addr, prefix, prefix_len, action_id, egress_p);
    endtask

    // ==========================================
    // Task: Send IPv4 packet with specified protocol
    // ==========================================
    task send_ipv4_packet(
        input [47:0] dst_mac,
        input [47:0] src_mac,
        input [31:0] src_ip,
        input [31:0] dst_ip,
        input [7:0]  protocol,
        input [7:0]  ttl,
        input [5:0]  dscp_in,
        input string description
    );
        logic [DATA_WIDTH-1:0] packet;

        packet = '0;

        // Ethernet header (14 bytes) - same format as working basic testbench
        packet[47:0]    = dst_mac;
        packet[95:48]   = src_mac;
        packet[111:96]  = 16'h0800;   // EtherType IPv4

        // IPv4 header (20 bytes) starting at byte 14
        // Byte 14: {IHL[3:0], Version[3:0]} = bits [119:112]
        // Byte 15: {DSCP[5:0], ECN[1:0]} = bits [127:120]
        packet[115:112] = 4'd4;       // version
        packet[119:116] = 4'd5;       // ihl
        packet[127:122] = dscp_in;    // DSCP (diffserv) - upper 6 bits of TOS
        packet[121:120] = 2'b00;      // ECN - lower 2 bits of TOS
        packet[143:128] = 16'd40;     // total length
        packet[159:144] = 16'h0001;   // identification
        packet[175:160] = 16'h4000;   // flags + frag offset (DF bit set)
        packet[183:176] = ttl;        // TTL
        packet[191:184] = protocol;   // protocol
        packet[207:192] = 16'h0000;   // checksum (placeholder)
        packet[239:208] = src_ip;     // src IP (wire order - same as basic)
        packet[271:240] = dst_ip;     // dst IP (wire order - same as basic)

        // Add L4 header placeholder
        if (protocol == PROTO_UDP) begin
            packet[287:272] = 16'd1234;   // src port
            packet[303:288] = 16'd5678;   // dst port
            packet[319:304] = 16'd20;     // length
            packet[335:320] = 16'd0;      // checksum
        end else if (protocol == PROTO_TCP) begin
            packet[287:272] = 16'd1234;   // src port
            packet[303:288] = 16'd80;     // dst port
            packet[335:304] = 32'h0;      // seq
            packet[367:336] = 32'h0;      // ack
            packet[375:368] = 8'h50;      // data offset + reserved
            packet[383:376] = 8'h02;      // flags (SYN)
        end

        ingress_port <= 9'd0;

        @(posedge aclk);
        s_axis_tvalid <= 1'b1;
        s_axis_tdata  <= packet;
        s_axis_tkeep  <= {KEEP_WIDTH{1'b1}};
        s_axis_tlast  <= 1'b1;

        wait(s_axis_tready);
        @(posedge aclk);
        s_axis_tvalid <= 1'b0;
        s_axis_tlast  <= 1'b0;

        packets_sent++;
        $display("[%0t] Sent packet #%0d: %s", $time, packets_sent, description);
        $display("        proto=%0d dscp_in=%0d dst_ip=%08h", protocol, dscp_in, dst_ip);
    endtask

    // ==========================================
    // Output monitor - check DSCP values
    // ==========================================
    always @(posedge aclk) begin
        if (m_axis_tvalid && m_axis_tready && m_axis_tlast) begin
            automatic logic [5:0] recv_dscp;
            automatic logic [7:0] recv_proto;

            // Extract DSCP from IPv4 header TOS byte (byte 15)
            // TOS byte layout: {DSCP[5:0], ECN[1:0]} at bits [127:120]
            // DSCP is upper 6 bits: [127:122]
            recv_dscp = m_axis_tdata[127:122];
            recv_proto = m_axis_tdata[191:184];

            packets_received++;
            $display("[%0t] Received packet #%0d:", $time, packets_received);
            $display("        Protocol: %0d, Output DSCP: %0d", recv_proto, recv_dscp);

            // Verify expected DSCP values
            if (recv_proto == PROTO_UDP && recv_dscp != DSCP_EF) begin
                $display("        WARNING: UDP should have DSCP=%0d (EF), got %0d", DSCP_EF, recv_dscp);
            end
            if (recv_proto == PROTO_TCP && recv_dscp != DSCP_VA) begin
                $display("        WARNING: TCP should have DSCP=%0d (VA), got %0d", DSCP_VA, recv_dscp);
            end
        end
    end

    // ==========================================
    // Debug: Parser outputs
    // ==========================================
    always @(posedge aclk) begin
        if (parser_payload_valid) begin
            $display("[%0t] PARSER: ipv4_valid=%b protocol=%0d dscp=%0d",
                    $time, ipv4_valid, ipv4_protocol, ipv4_diffserv);
        end
    end

    // ==========================================
    // Debug: QoS DSCP marking
    // ==========================================
    always @(posedge aclk) begin
        if (match_action_inst.match_valid) begin
            $display("[%0t] MATCH-ACTION: action=%0d qos_udp=%b qos_tcp=%b dscp_out=%0d",
                    $time,
                    match_action_inst.match_action_id,
                    match_action_inst.qos_cond_1_match,  // UDP condition
                    match_action_inst.qos_cond_2_match,  // TCP condition
                    pipeline_ipv4_diffserv);
        end
    end

    // ==========================================
    // Main test sequence
    // ==========================================
    initial begin
        // Initialize signals
        s_axis_tvalid = 0;
        s_axis_tdata  = 0;
        s_axis_tkeep  = 0;
        s_axis_tlast  = 0;
        m_axis_tready = 1;
        table_wr_en   = 0;
        table_wr_addr = 0;
        table_entry_valid = 0;
        table_entry_prefix = 0;
        table_entry_prefix_len = 0;
        table_entry_action = 0;
        table_entry_action_data = 0;
        ingress_port  = 9'd0;

        // Wait for reset release
        @(posedge aresetn);
        repeat(10) @(posedge aclk);

        $display("\n========================================================");
        $display("           QoS (DSCP Marking) Testbench");
        $display("========================================================");
        $display("Expected QoS marking behavior:");
        $display("  - UDP packets (proto=17) -> DSCP=%0d (Expedited Forwarding)", DSCP_EF);
        $display("  - TCP packets (proto=6)  -> DSCP=%0d (Voice Admit)", DSCP_VA);
        $display("  - Other protocols        -> DSCP unchanged");
        $display("========================================================\n");

        // ========================================
        // Configure routing table
        // IP prefixes in BIG-ENDIAN (network order) to match parser output
        // ========================================
        $display("Configuring routing table...\n");

        // Route for 10.0.0.0/8 -> forward to port 1
        configure_route(
            .addr(0),
            .prefix(32'h0A000000),  // 10.0.0.0 in big-endian (network order)
            .prefix_len(6'd8),
            .action_id(ACTION_FORWARD),
            .dst_mac(48'hAABBCCDDEE01),
            .egress_p(9'd1)
        );

        // Route for 192.168.1.0/24 -> forward to port 2
        configure_route(
            .addr(1),
            .prefix(32'hC0A80100),  // 192.168.1.0 in big-endian (network order)
            .prefix_len(6'd24),
            .action_id(ACTION_FORWARD),
            .dst_mac(48'hAABBCCDDEE02),
            .egress_p(9'd2)
        );

        repeat(10) @(posedge aclk);

        // ========================================
        // Test Cases
        // ========================================

        // Test 1: UDP packet -> should get DSCP=46 (Expedited Forwarding)
        $display("\n--- Test 1: UDP packet -> DSCP=46 (EF) ---");
        send_ipv4_packet(
            .dst_mac(48'hFFFFFFFFFFFF),
            .src_mac(48'h112233445566),
            .src_ip(32'h0101A8C0),    // 192.168.1.1 (little-endian, parser will bswap)
            .dst_ip(32'h0100000A),    // 10.0.0.1 (little-endian)
            .protocol(PROTO_UDP),
            .ttl(8'd64),
            .dscp_in(6'd0),
            .description("UDP packet to 10.0.0.1")
        );
        repeat(30) @(posedge aclk);

        // Test 2: TCP packet -> should get DSCP=44 (Voice Admit)
        $display("\n--- Test 2: TCP packet -> DSCP=44 (VA) ---");
        send_ipv4_packet(
            .dst_mac(48'hFFFFFFFFFFFF),
            .src_mac(48'h112233445566),
            .src_ip(32'h0201A8C0),    // 192.168.1.2 (little-endian)
            .dst_ip(32'h0200000A),    // 10.0.0.2 (little-endian)
            .protocol(PROTO_TCP),
            .ttl(8'd64),
            .dscp_in(6'd0),
            .description("TCP packet to 10.0.0.2")
        );
        repeat(30) @(posedge aclk);

        // Test 3: ICMP packet -> DSCP should remain 0 (no QoS marking)
        $display("\n--- Test 3: ICMP packet -> DSCP unchanged (0) ---");
        send_ipv4_packet(
            .dst_mac(48'hFFFFFFFFFFFF),
            .src_mac(48'h112233445566),
            .src_ip(32'h0301A8C0),    // 192.168.1.3 (little-endian)
            .dst_ip(32'h0300000A),    // 10.0.0.3 (little-endian)
            .protocol(PROTO_ICMP),
            .ttl(8'd64),
            .dscp_in(6'd0),
            .description("ICMP packet to 10.0.0.3")
        );
        repeat(30) @(posedge aclk);

        // Test 4: UDP packet with existing DSCP -> should override to 46
        $display("\n--- Test 4: UDP with DSCP=10 -> should override to DSCP=46 ---");
        send_ipv4_packet(
            .dst_mac(48'hFFFFFFFFFFFF),
            .src_mac(48'h112233445566),
            .src_ip(32'h0401A8C0),    // 192.168.1.4 (little-endian)
            .dst_ip(32'h6401A8C0),    // 192.168.1.100 (little-endian)
            .protocol(PROTO_UDP),
            .ttl(8'd64),
            .dscp_in(6'd10),          // AF11 - should be overwritten
            .description("UDP with pre-set DSCP=10")
        );
        repeat(30) @(posedge aclk);

        // Test 5: TCP packet to different destination
        $display("\n--- Test 5: TCP to 192.168.1.x network -> DSCP=44 ---");
        send_ipv4_packet(
            .dst_mac(48'hFFFFFFFFFFFF),
            .src_mac(48'h112233445566),
            .src_ip(32'h0100000A),    // 10.0.0.1 (little-endian)
            .dst_ip(32'h0501A8C0),    // 192.168.1.5 (little-endian)
            .protocol(PROTO_TCP),
            .ttl(8'd64),
            .dscp_in(6'd0),
            .description("TCP packet to 192.168.1.5")
        );
        repeat(30) @(posedge aclk);

        // Test 6: UDP with high DSCP -> should still override
        $display("\n--- Test 6: UDP with DSCP=46 (already EF) -> remains 46 ---");
        send_ipv4_packet(
            .dst_mac(48'hFFFFFFFFFFFF),
            .src_mac(48'h112233445566),
            .src_ip(32'h0601A8C0),    // 192.168.1.6 (little-endian)
            .dst_ip(32'h0600000A),    // 10.0.0.6 (little-endian)
            .protocol(PROTO_UDP),
            .ttl(8'd64),
            .dscp_in(6'd46),
            .description("UDP with pre-set DSCP=46")
        );
        repeat(30) @(posedge aclk);

        // ========================================
        // Final Summary
        // ========================================
        repeat(50) @(posedge aclk);

        $display("\n========================================================");
        $display("                    Test Summary");
        $display("========================================================");
        $display("Packets sent:     %0d", packets_sent);
        $display("Packets received: %0d", packets_received);
        $display("Total processed:  %0d", packet_count);
        $display("Forwarded:        %0d", forwarded_count);
        $display("Dropped:          %0d", dropped_count);
        $display("========================================================");
        $display("\nExpected Results:");
        $display("  - Test 1 (UDP):  DSCP=46 (Expedited Forwarding)");
        $display("  - Test 2 (TCP):  DSCP=44 (Voice Admit)");
        $display("  - Test 3 (ICMP): DSCP=0 (unchanged)");
        $display("  - Test 4 (UDP):  DSCP=46 (override from 10)");
        $display("  - Test 5 (TCP):  DSCP=44 (Voice Admit)");
        $display("  - Test 6 (UDP):  DSCP=46 (remains 46)");
        $display("========================================================\n");

        if (packets_received == packets_sent && packets_sent > 0) begin
            $display("*** TEST PASSED ***\n");
        end else begin
            $display("*** TEST FAILED ***\n");
        end

        $finish;
    end

endmodule
